module lowpass(
    input wire clk,
    input wire rst,
    input wire signed
)

